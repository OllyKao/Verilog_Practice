module top_module (
    input clk,
    input reset,            // Synchronous reset
    input [7:0] d,
    output [7:0] q
);

    always @(posedge clk) begin
        q <= (reset == 1'b1)? 7'b0 : d;
    end

endmodule

module top_module(
    input clk,
    input [7:0] in,
    input reset,    // Synchronous reset
    output [23:0] out_bytes,
    output done); //
    
	reg [1:0] state, next_state;
    
    // FSM from fsm_ps2
    always @(*) begin
        case(state)
            2'b00:	next_state = in[3]? 2'b01 : 2'b00;
            2'b01:	next_state = 2'b10;
            2'b10:	next_state = 2'b11;
            2'b11:	next_state = in[3]? 2'b01 : 2'b00;
        endcase
    end
   
    always @(posedge clk) begin
        if(reset)
            state <= 2'b0;
        else begin
            state <= next_state;
            out_bytes[((4 - next_state) * 8 - 1) -:8] <= in;
        end
    end
 
    assign done = (state == 2'b11);

endmodule
